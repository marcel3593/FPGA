`define EEPROM_NOP      2'b00
`define EEPROM_WR       2'b01
`define EEPROM_RD       2'b10
`define EEPROM_LDA      2'b11