    .INIT_00(256'h0000002fb1809c0800000006b2009d080000000b21809e0800000014b0009f08),
    .INIT_01(256'h00000020a5500ce00000000b92d2063b0000000b82c00cd0000000001502063b),
    .INIT_02(256'h0000000ba252066100000001b002063b00000020a7f00cf000000020a612063b),
    .INIT_03(256'h00000014a00224920000000ba262085e00000014b003640000000014a0e19201),
    .INIT_04(256'h00000014a00206b800000014b002069f00000014a003649300000014b001d050),
    .INIT_05(256'h0000002f21b20663000000062b0364910000000b21b1d02000000014b0009006),
    .INIT_06(256'h00000014b002062000000014a003a49100000014b002065100000014a0001202),
    .INIT_07(256'h00000014b002062000000014a002fb1300000014b002062000000014a0020620),
    .INIT_08(256'h00000014a00364590000000ba270d04000000014b000900200000014a0020620),
    .INIT_09(256'h00000014a003245900000014b001fb0000000014a001da0000000014b0003b03),
    .INIT_0A(256'h0000002fb1a1da8000000006b20324590000000b21a1fb0000000014b001da20),
    .INIT_0B(256'h00000020a551fb000000000b92f1daa00000000b82e32459000000001401fb00),
    .INIT_0C(256'h0000000ba253245900000001b001fb0000000020a7f1dac000000020a6132459),
    .INIT_0D(256'h00000014a001da200000000ba263245900000014b001fb0000000014a0e1dae0),
    .INIT_0E(256'h00000014a001fb0100000014b001da8000000014a003245900000014b001fb01),
    .INIT_0F(256'h0000002f21d32459000000062b01fb010000000b21d1daa000000014b0032459),
    .INIT_10(256'h00000014b001da0000000014a003245900000014b001fb0100000014a001dac0),
    .INIT_11(256'h00000014b001fb0200000014a001da2000000014b003245900000014a001fb02),
    .INIT_12(256'h00000014a00324590000000ba271fb0200000014b001da8000000014a0032459),
    .INIT_13(256'h00000014a001dac000000014b003245900000014a001fb0200000014b001daa0),
    .INIT_14(256'h0000002fb1c1fb0300000006b201da000000000b21c3245900000014b001fb02),
    .INIT_15(256'h0000000d1ff3245900000001b001fb0300000001a001dae00000002500032459),
    .INIT_16(256'h0000000d9ff0b01300000014a002088a0000000d8ff2066100000014a0022491),
    .INIT_17(256'h0000002fb253246900000014b001d0010000000daff3246400000014a001d000),
    .INIT_18(256'h0000000d1ff3247b00000001a001d0030000000020032471000000250001d002),
    .INIT_19(256'h00000014a04208e500000014a04208ba00000014a04001b000000014a00000a0),
    .INIT_1A(256'h00000014a04207a200000014a042085800000014a04207a200000014a0422486),
    .INIT_1B(256'h000000062b0208e500000020a72208ba000000022a0001b000000014a04000a0),
    .INIT_1C(256'h00000000b90207a200000000a802085800000025000207a20000002f22622486),
    .INIT_1D(256'h00000014b00001b000000014a06000a000000014b00207a200000014a0620858),
    .INIT_1E(256'h00000014b00207a200000014a062248600000014b00208e500000014a06208ba),
    .INIT_1F(256'h00000000210207a2000000250002085800000014b00207a200000014a0620858),
    .INIT_20(256'h000000032aa001b000000001b00000a000000001a00207a20000000038020858),
    .INIT_21(256'h0000000d3ff00cf000000014a0000bc00000000d2ff208e500000003301208ba),
    .INIT_22(256'h0000000021000cd000000014b082063b0000000daff00ce000000014a002063b),
    .INIT_23(256'h000000033022085e000000032cc2063b00000001a0000cb0000000003802063b),
    .INIT_24(256'h00000014a002200a0000000d3ff2071600000014a00206610000000d2ff22491),
    .INIT_25(256'h0000000038020076000000002102006d00000014b08206610000000daff2069d),
    .INIT_26(256'h0000000d2ff2007f00000003304324a0000000032f01d00200000001a000b002),
    .INIT_27(256'h0000000daff2008800000014a00324a00000000d3ff1d00300000014a000b002),
    .INIT_28(256'h000000370012071600000025000206d50000002fb270100200000014b082085e),
    .INIT_29(256'h0000000b40e200760000000b30d2006d0000000b20c2066100000020b912200a),
    .INIT_2A(256'h0000001450e2007f00000003403324b0000000005401d0020000000ba0f0b002),
    .INIT_2B(256'h000000007a02008800000003607324b0000000006a01d0030000001450e0b002),
    .INIT_2C(256'h0000001470e010010000001470e2f01e0000001470e010000000001470e2085e),
    .INIT_2D(256'h000000008202066700000001e002068700000001d00206f1000000037032f032),
    .INIT_2E(256'h00000032b072088a0000001d6032066100000032adf225440000001d60220663),
    .INIT_2F(256'h00000001a002259100000001900206f100000032b472f0320000001d60401002),
    .INIT_30(256'h00000032acb206420000001ce400bc3300000036ac4206630000001cd302069b),
    .INIT_31(256'h00000013a000bc0b00000013900206b5000000108f02064c00000009f0820642),
    .INIT_32(256'h00000001d000bc0900000022ac02063b00000013e000bc0a00000011d012063b),
    .INIT_33(256'h00000032ad50bc070000001cd502063b0000000bf310bc080000000be302063b),
    .INIT_34(256'h00000011d010d00800000013a0009002000000129f020661000000108e02063b),
    .INIT_35(256'h00000003a03206d50000002f911010100000002f8102088a00000022ace324d9),
    .INIT_36(256'h00000004a002071600000014006206d500000014006010000000000b0132200a),
    .INIT_37(256'h0000000bd300bc09000000250000bb08000000370000ba070000002fa122200a),
    .INIT_38(256'h00000001a00000f0000000019000bf330000000b2370be0b0000000be310bd0a),
    .INIT_39(256'h000000108d00d00800000032aec324ea0000001cf201d00c00000001f000300f),
    .INIT_3A(256'h00000022ae50301f00000011f01000a000000013a002253f000000129e0324ea),
    .INIT_3B(256'h00000032af5206200000001cf50206200000000b23c2062000000001f002f014),
    .INIT_3C(256'h00000011f013e53f00000013a001d05d000000139000307f00000010820000b0),
    .INIT_3D(256'h00000032afd1d00c0000001cf300300f00000001f000b03300000022aee2f015),
    .INIT_3E(256'h00000011f01000e00000001380032504000000139000d00800000011802324fb),
    .INIT_3F(256'h00000003a030b1130000002f9112f0130000002f8100300300000022af61400e),
    .INIT_40(256'h00000004a00365130000001400620620000000140063653f0000000b0131c010),
    .INIT_41(256'h0000000bd300b113000000250002f01300000037000030030000002fa120b033),
    .INIT_42(256'h000000019002fc0c00000001800206200000000b2373653f0000000be311c010),
    .INIT_43(256'h00000032b1503f070000001cf202ff0f00000001f002fe0e00000001a002fd0d),
    .INIT_44(256'h00000011f0103e0300000013a0022523000000129e03253f000000108d01df01),
    .INIT_45(256'h0000001df0020b9100000003ff02fe120000000bf392fd1100000022b0e2fc10),
    .INIT_46(256'h0000000b01318c000000000b23c0b20600000001f000b10500000032b2c0b004),
    .INIT_47(256'h00000032b2c20bbc0000001df023e53f00000032b251ae200000001d0001ad10),
    .INIT_48(256'h00000011f010b01300000013a002f40f0000001390003407000000108200b40f),
    .INIT_49(256'h000000108203253100000032b2c1d0010000001df013252c00000022b1e1d000),
    .INIT_4A(256'h00000022b253253b00000011f011d00300000013a0032536000000139001d002),
    .INIT_4B(256'h00000032b35209000000001cf50206050000000b238207d000000001f00208eb),
    .INIT_4C(256'h00000011f012060500000013a00207d700000013900208ee000000108202253f),
    .INIT_4D(256'h00000032b3d207e10000001cf30208f100000001f002253f00000022b2e2090a),
    .INIT_4E(256'h00000011f01208f4000000138002253f00000013900209150000001180120605),
    .INIT_4F(256'h00000003a032085e0000002f911209200000002f8102060500000022b36207ed),
    .INIT_50(256'h00000004a002200a000000140062071600000014006206d50000000b01301000),
    .INIT_51(256'h0000000bd300900e0000002500036097000000370000d0080000002fa1209011),
    .INIT_52(256'h0000000190036103000000018000d0400000000b237361070000000be310d080),
    .INIT_53(256'h00000032b55360fb0000001cf200d01000000001f00360ff00000001a000d020),
    .INIT_54(256'h00000011f010901600000013a003255a000000129e00d004000000108d00900e),
    .INIT_55(256'h0000001df001d00e00000003ff00300f0000000bf392b04e00000022b4e2f033),
    .INIT_56(256'h0000000b0130d0200000000b23c0900d00000001f002254400000032b6c3256e),
    .INIT_57(256'h00000032b6c3256e0000001df021d04900000032b65090060000001d00036544),
    .INIT_58(256'h00000011f012066100000013a00206a50000001390036544000000108201d053),
    .INIT_59(256'h000000108201130100000032b6c2071f0000001df010130000000022b5e0b202),
    .INIT_5A(256'h00000022b652066700000011f012068700000013a0036566000000139001c320),
    .INIT_5B(256'h0000001cf00206610000000b037206910000000b2382254400000001f0020663),
    .INIT_5C(256'h00000013a001d002000000139000b002000000108202004700000032b762003e),
    .INIT_5D(256'h0000000b2031d00300000001f000b00200000022b6e2005000000011f013257a),
    .INIT_5E(256'h0000001390022589000000108202085e00000032b7f200590000001cf503257a),
    .INIT_5F(256'h00000001f001d00200000022b780b00200000011f012004700000013a002003e),
    .INIT_60(256'h000000139001d003000000118010b00200000032b87200500000001cf3032586),
    .INIT_61(256'h0000002f8100106000000022b802085e00000011f01200590000001380032586),
    .INIT_62(256'h000000140062d0030000000b0132f03200000003a03010000000002f911206c9),
    .INIT_63(256'h00000037000207160000002fa12206d500000004a00010000000001400620703),
    .INIT_64(256'h00000032b9801f000000001d00001e000000000b01301d00000000250002200a),
    .INIT_65(256'h00000032b9a01d000000001d0302ff12000000030f02fe110000000b0392fd10),
    .INIT_66(256'h000000095082fd1e00000020bb501d0100000022b9b2fd1300000020bae2fd01),
    .INIT_67(256'h0000002f504325bc000000096081d0ff000000095080b00f0000002f50320bbc),
    .INIT_68(256'h0000002f5300b001000000096082f00f00000009508030070000002f6050b00f),
    .INIT_69(256'h0000002f537325b0000000096081d00100000009508325ac0000002f6311d000),
    .INIT_6A(256'h0000002f53c325b8000000096081d00300000009508325b40000002f6381d002),
    .INIT_6B(256'h0000000160722172000000015ef2093f00000025000207d00000002f606208eb),
    .INIT_6C(256'h0000002d10b221720000002d60a2093f0000002d509207d700000001100208ee),
    .INIT_6D(256'h00000001100221720000000160b2093f000000015c3207e100000025000208f1),
    .INIT_6E(256'h00000025000221720000002d10b2093f0000002d60a207ed0000002d509208f4),
    .INIT_6F(256'h0000000b911090160000000b810325c500000020b910d004000000370010900e),
    .INIT_70(256'h0000002fa361d00e0000002f9350300f0000002f8342b04e0000000ba122f033),
    .INIT_71(256'h0000000b4310b1050000000b3300b0040000000bd3720b9100000001200325e7),
    .INIT_72(256'h0000003abd30bf120000001ba000be110000001a9400bd10000000188300b206),
    .INIT_73(256'h0000002fa361ef200000002f9351ee100000002f8341cd000000001120103f03),
    .INIT_74(256'h0000000b83413f0000000022bc813e0000000032bff11d010000001c2d0325d8),
    .INIT_75(256'h000000012002259a0000002f20f2ff120000000ba362fe110000000b9352fd10),
    .INIT_76(256'h00000032c971c0100000001d40119101000000094080b102000000013000b001),
    .INIT_77(256'h0000003abe62f0130000001ba002f0010000001b9001100100000018840325e7),
    .INIT_78(256'h0000002f9352fd100000002f83401f000000001330001e000000001120101d00),
    .INIT_79(256'h0000000b935207a20000000b8342259a00000022bd92ff120000002fa362fe11),
    .INIT_7A(256'h0000002f80c2d0030000002f20d010000000002f30e207b20000000ba3620037),
    .INIT_7B(256'h0000000b70f2200a0000000b60e207160000000b50d206d50000000b40c01000),
    .INIT_7C(256'h000000147002500000000014608365f0000000146080d0800000000b30e0900d),
    .INIT_7D(256'h0000000b013250000000002f70e365f4000000147000d040000000143080900d),
    .INIT_7E(256'h000000140062de0700000014006205f4000000140062df0700000014006205f4),
    .INIT_7F(256'h0000000b4392dc0700000025000205f4000000370002dd070000002f00f205f4),
    .INITP_00(256'hbf8abf9cbf8e341997098ca79eb78aa48bbfaa06aa12141e84b08d081cac12be),
    .INITP_01(256'h9a01183807351b241024a78da582931113a31d060f249d331ba79a368f3d219c),
    .INITP_02(256'h80a5be053808148d1e84b2b91ca585221d3801bf1b24351b22103801b91b241d),
    .INITP_03(256'ha221bb04bb032d8ca181bb0405a33a98081e331a849f849812179e0611263222),
    .INITP_04(256'hb81ba2119a8fa934b92eaab50630140f933db4312aaab7143b158c999200bda6),
    .INITP_05(256'ha5b3a3851b1bbb842e1a963d2b20a8ba03813f8f863927b6862d14ad2abf143e),
    .INITP_06(256'h8aa32aa13a18973c11ba9088222490853ca3b71789110b22ad3d930c2a210a1b),
    .INITP_07(256'h1ab91f859f14b52930abb21b87a3af1db58f1dbb9394a48804a2b725a12e181c),
    .INITP_08(256'h1b051d852718bf020882293f05ac8e8b0a3ea0a3aa1d9d0792ba2636a0990524),
    .INITP_09(256'h8c208b379600262301aca1a981b3ae10020088292e91362102968aa489b92f0e),
    .INITP_0A(256'h249ab206a304a8248a0fab0c9f368f9334a926bcaf9916860721b52aad9418a8),
    .INITP_0B(256'ha3898eb6af123f8903329408a6b08eb938a916b28a8820bf96a4001f8633a813),
    .INITP_0C(256'h249705ac1faa0e2d3508002ea08dbba430ba3918872b9eb48b07031da221a432),
    .INITP_0D(256'ha90f3e38a6381b0d80b5b6a3b3809c8bbf32b72cbe920f3da517813fb08117b4),
    .INITP_0E(256'h27188c9b932f293782022caa143c1888b7bf1f283d8283bf07319a9ea5a49730),
    .INITP_0F(256'h1cb5b63711121c12ab1e381db19e013d812fa513058dacb53f1fb929af14a133),
